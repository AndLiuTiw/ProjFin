// NOTE : Below mentioned frame work is for reference purpose.
module simplified_sha256 #(parameter integer NUM_OF_WORDS = 20)(
 input logic  clk, reset_n, start,
 input logic  [15:0] message_addr, output_addr,
 output logic done, mem_clk, mem_we,
 output logic [15:0] mem_addr,
 output logic [31:0] mem_write_data,
 input logic [31:0] mem_read_data);

// FSM state variables 
enum logic [2:0] {IDLE, READ, BLOCK, COMPUTE, WRITE} state;
enum logic [1:0] {EXPAND, OP, OUT} step;

// NOTE : Below mentioned frame work is for reference purpose.
// Local variables might not be complete and you might have to add more variables
// or modify these variables. Code below is more as a reference.

// Local variables
logic [31:0] w[16]; //To be used in word expansion and sha operation steps, have not initialized yet
logic [31:0] message[20]; //These are the 20 message blocks, each one is 32 bits
logic [31:0] wt; //Wtf is this (unused for now)
logic [31:0] h0, h1, h2, h3, h4, h5, h6, h7; //initialized in always_ff block BLOCK state
logic [31:0] a, b, c, d, e, f, g, h; //initialized in always_ff block IDLE state
logic [ 7:0] i, j, ind, ind2; //i has been initialized in IDLE, we're using j as the index variable to load different blocks, ind is being used in the WRITE state, ind2 is being usd in the READ state
logic [15:0] offset; // in word address //initialized in IDLE state
logic        cur_we; //initialized in IDLE state 
logic [15:0] cur_addr; //Initialized in IDLE state
logic [31:0] cur_write_data; //Unitialized, it's use is understood
logic [511:0] memory_block; //Not sure how this is to be used (unitialized)

// SHA256 K constants
parameter int k[0:63] = '{
   32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
   32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
   32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
   32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
   32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
   32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
   32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
   32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};


// Generate request to memory
// for reading from memory to get original message
// for writing final computed has value
assign mem_clk = clk;
assign mem_addr = cur_addr + offset; 
assign mem_we = cur_we;
assign mem_write_data = cur_write_data;


// Right Rotation Example : right rotate input x by r
// Lets say input x = 1111 ffff 2222 3333 4444 6666 7777 8888
// lets say r = 4
// x >> r  will result in : 0000 1111 ffff 2222 3333 4444 6666 7777 
// x << (32-r) will result in : 8888 0000 0000 0000 0000 0000 0000 0000
// final right rotate expression is = (x >> r) | (x << (32-r));
// (0000 1111 ffff 2222 3333 4444 6666 7777) | (8888 0000 0000 0000 0000 0000 0000 0000)
// final value after right rotate = 8888 1111 ffff 2222 3333 4444 6666 7777
// Right rotation function
function logic [31:0] rightrotate(input logic [31:0] x,
                                  input logic [ 7:0] r);
   rightrotate = (x >> r) | (x << (32 - r));
endfunction


// SHA-256 FSM 
// Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
// and write back hash value back to memory
always_ff @(posedge clk, negedge reset_n)
begin
  if (!reset_n) begin
    cur_we <= 1'b0;
    state <= IDLE;
  end 
  else case (state)
    // Initialize hash values h0 to h7 and a to h, other variables and memory we, address offset, etc
    IDLE: begin 
       if(start) begin
       // Student to add rest of the code
		   //a through h are initialized to initial hash values
			a <= 32'h6a09e667; 
			b <= 32'hbb67ae85;
			c <= 32'h3c6ef372;
			d <= 32'ha54ff53a;
			e <= 32'h510e527f;
			f <= 32'h9b05688c;
			g <= 32'h1f83d9ab;
			h <= 32'h5be0cd19;
			cur_we <= 0; //Because nothing needs to be written to memory right now (in the idle state)
			offset <= 0; //Should probably be 0 initially
			cur_addr <= message_addr; //Because curr_addr should be initialized to 1st message location (address of W0 (We have words from W0 to W15))in memory
			j <= 0; //used
			ind2 <= 0; //Because next state is the READ state
			offset <= 0; //Because next state is READ state and I need to create a 1 cycle gap
			state <= READ;
       end
    end
	 
	 //Adding a READ state to Read 640 bits message from testbench memory in chunks of 32bits words (i.e. read 20 locations from memory by incrementing address offset)
	 READ: begin
		if(ind2 > 0) begin
			message[ind2 - 1] <= mem_read_data;
		end
		if(ind2 <= 19) begin
			offset <= offset + 16'd1; //To read from next address in memory
			ind2 <= ind2 + 8'd1;
			state <= READ;
		end
		else begin
			state <= BLOCK;
		end
	 end

    // SHA-256 FSM 
    // Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function    
    // and write back hash value back to memory
    BLOCK: begin
	// Fetch message in 512-bit block size
	// For each of 512-bit block initiate hash value computation
	   h0 <= a;
		h1 <= b;
		h2 <= c;
		h3 <= d;
		h4 <= e;
		h5 <= f;
		h6 <= g;
		h7 <= h;
		if (j == 0) begin 
			for (int n = 0; n < 16; n++) begin
				w[n] <= message[n];
			end
			j <= j + 8'd1;
			state <= COMPUTE;
			i <= 0;
			step <= OP;
		end
		else if (j == 1) begin
			for (int n = 0; n < 4; n++) begin
				w[n] <= message[n+16];
			end
			w[4] <= 32'h80000000;
			for (int n = 0; n < 10; n++) begin
				w[n+5] <= 32'b0;
			end
			w[15] <= 32'd640;
			j <= j + 8'd1;
			state <= COMPUTE;
			i <= 0;
			step <= OP;
		end
		else if(j == 2) begin //This is to create a 1 cycle delay so that the right value of h0 can be written
			j <=  j + 8'd1;
			state <= BLOCK;
		end
		else begin //j is equal to 3
			cur_we <= 1; //Because the next state is the WRITE state
			cur_addr <= output_addr; //Because the next state is the WRITE state
			offset <= 0; //Because the next state is the WRITE state
			ind <= 0; //Because the next state is the WRITE state
			cur_write_data <= h0; //Will be written at next clock edge
			state <= WRITE;
		end
    end

    // For each block compute hash function
    // Go back to BLOCK stage after each block hash computation is completed and if
    // there are still number of message blocks available in memory otherwise
    // move to WRITE stage
	COMPUTE: begin
	// 64 processing rounds steps for 512-bit block
		// shift w every time to keep the useful 16 words in it
		case(step)
			OP: begin
			// this is the word expansion part
				// store w_new at w 
				for (int n = 0; n < 15; n++) begin
					w[n] <= w[n+1];
				end
				w[15] <= w[0] 
					+ w[9]
					+ (rightrotate(w[1],7) ^ rightrotate(w[1],18) ^ (w[1] >> 3)) 
					+ (rightrotate(w[14],17) ^ rightrotate(w[14],19) ^ (w[14] >> 10));
//				w[15] <= wt;
			// this is the sha256_op part
				a <= h 
					+ (rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25)) 
					+ ((e & f) ^ ((~e) & g)) + k[i] + w[0] 
					+ (rightrotate(a, 2) ^ rightrotate(a, 13) ^ rightrotate(a, 22)) 
					+ ((a & b) ^ (a & c) ^ (b & c));
				b <= a;
				c <= b;
				d <= c;
				e <= d 
					+ h 
					+ (rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25)) 
					+ ((e & f) ^ ((~e) & g)) 
					+ k[i] 
					+ w[0];
				f <= e;
				g <= f;
				h <= g;
				i <= i + 8'd1;
				if (i == 63) begin
					step <= OUT;
				end
				state <= COMPUTE; //Go back to compute if i value is in [65, 128]
			end
			OUT: begin
			// for last compression
				//a through h are going to be used again BLOCK state to initialize h0 to h7
				a <= a + h0;
				b <= b + h1;
				c <= c + h2;
				d <= d + h3;
				e <= e + h4;
				f <= f + h5;
				g <= g + h6;
				h <= h + h7;
				state <= BLOCK; //Go to BLOCK state if i value is 129
			end
		endcase
	end

    // h0 to h7 each are 32 bit hashes, which makes up total 256 bit value
    // h0 to h7 after compute stage has final computed hash value
    // write back these h0 to h7 to memory starting from output_addr
    WRITE: begin
		case (ind)
			0 : begin
				offset <= 1;
				cur_write_data <= h1;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			1 : begin
				offset <= 2;
				cur_write_data <= h2;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			2 : begin
				offset <= 3;
				cur_write_data <= h3;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			3 : begin
				offset <= 4;
				cur_write_data <= h4;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			4 : begin
				offset <= 5;
				cur_write_data <= h5;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			5 : begin
				offset <= 6;
				cur_write_data <= h6;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			6 : begin
				offset <= 7;
				cur_write_data <= h7;
				ind <= ind + 8'd1;
				state <= WRITE;
			end
			7 : begin
				offset <= 0;
				cur_we <= 0; //Because next state is IDLE state
				ind <= 8'd0;
				state <= IDLE;
			end
		endcase
    end
   endcase
  end

//assign sha256_func_output = sha256_op(a, b, c, d, e, f, g, h, w, tstep);
// Generate done when SHA256 hash computation has finished and moved to IDLE state
assign done = (state == IDLE);

endmodule
